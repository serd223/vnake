module snake

pub enum Direction {
	up
	down
	left
	right
	stopped
}
